
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hd57c2016;
    ram_cell[       1] = 32'h0;  // 32'h661f505a;
    ram_cell[       2] = 32'h0;  // 32'h71eef11e;
    ram_cell[       3] = 32'h0;  // 32'hb852580e;
    ram_cell[       4] = 32'h0;  // 32'h79a29c4d;
    ram_cell[       5] = 32'h0;  // 32'hea6ceefa;
    ram_cell[       6] = 32'h0;  // 32'hf9266cad;
    ram_cell[       7] = 32'h0;  // 32'h4dc699fb;
    ram_cell[       8] = 32'h0;  // 32'he777d506;
    ram_cell[       9] = 32'h0;  // 32'h45538379;
    ram_cell[      10] = 32'h0;  // 32'hd63a3016;
    ram_cell[      11] = 32'h0;  // 32'h6b4e7a47;
    ram_cell[      12] = 32'h0;  // 32'haa2fadd9;
    ram_cell[      13] = 32'h0;  // 32'h5660028f;
    ram_cell[      14] = 32'h0;  // 32'h61004602;
    ram_cell[      15] = 32'h0;  // 32'hc5263e95;
    ram_cell[      16] = 32'h0;  // 32'he7f1da1d;
    ram_cell[      17] = 32'h0;  // 32'ha51a38d4;
    ram_cell[      18] = 32'h0;  // 32'hfca4922c;
    ram_cell[      19] = 32'h0;  // 32'h33a0a6f8;
    ram_cell[      20] = 32'h0;  // 32'h6eb40359;
    ram_cell[      21] = 32'h0;  // 32'h0591d8cd;
    ram_cell[      22] = 32'h0;  // 32'he4385aaa;
    ram_cell[      23] = 32'h0;  // 32'hac7ce49e;
    ram_cell[      24] = 32'h0;  // 32'h113c5f24;
    ram_cell[      25] = 32'h0;  // 32'h29660181;
    ram_cell[      26] = 32'h0;  // 32'h706b7caf;
    ram_cell[      27] = 32'h0;  // 32'h5a46e192;
    ram_cell[      28] = 32'h0;  // 32'ha68bebef;
    ram_cell[      29] = 32'h0;  // 32'h45fa6851;
    ram_cell[      30] = 32'h0;  // 32'h06b6109a;
    ram_cell[      31] = 32'h0;  // 32'h6df0ad51;
    ram_cell[      32] = 32'h0;  // 32'h7a695799;
    ram_cell[      33] = 32'h0;  // 32'h72d28a34;
    ram_cell[      34] = 32'h0;  // 32'he8808334;
    ram_cell[      35] = 32'h0;  // 32'h9e1e1d8b;
    ram_cell[      36] = 32'h0;  // 32'hbe025244;
    ram_cell[      37] = 32'h0;  // 32'h29086f4f;
    ram_cell[      38] = 32'h0;  // 32'h2e8b2a2d;
    ram_cell[      39] = 32'h0;  // 32'h5e666470;
    ram_cell[      40] = 32'h0;  // 32'h1067676b;
    ram_cell[      41] = 32'h0;  // 32'hbd102e35;
    ram_cell[      42] = 32'h0;  // 32'hf3035e7a;
    ram_cell[      43] = 32'h0;  // 32'h31342d12;
    ram_cell[      44] = 32'h0;  // 32'h7e510fa5;
    ram_cell[      45] = 32'h0;  // 32'hadb37d92;
    ram_cell[      46] = 32'h0;  // 32'habde1992;
    ram_cell[      47] = 32'h0;  // 32'h378ce4bd;
    ram_cell[      48] = 32'h0;  // 32'h13b3a1be;
    ram_cell[      49] = 32'h0;  // 32'h037a7a5f;
    ram_cell[      50] = 32'h0;  // 32'hcc300bac;
    ram_cell[      51] = 32'h0;  // 32'h22c5cd43;
    ram_cell[      52] = 32'h0;  // 32'hedc69801;
    ram_cell[      53] = 32'h0;  // 32'hf46cf774;
    ram_cell[      54] = 32'h0;  // 32'ha8d6a585;
    ram_cell[      55] = 32'h0;  // 32'heee3499a;
    ram_cell[      56] = 32'h0;  // 32'he5466ab1;
    ram_cell[      57] = 32'h0;  // 32'h8fd52c91;
    ram_cell[      58] = 32'h0;  // 32'hcecdd7ee;
    ram_cell[      59] = 32'h0;  // 32'h3e0dee49;
    ram_cell[      60] = 32'h0;  // 32'h0efc6b3a;
    ram_cell[      61] = 32'h0;  // 32'he072596c;
    ram_cell[      62] = 32'h0;  // 32'h6e8493f2;
    ram_cell[      63] = 32'h0;  // 32'hc59fb143;
    ram_cell[      64] = 32'h0;  // 32'hbe2fd7e2;
    ram_cell[      65] = 32'h0;  // 32'ha3e9aeb7;
    ram_cell[      66] = 32'h0;  // 32'hd5c89963;
    ram_cell[      67] = 32'h0;  // 32'h2b999350;
    ram_cell[      68] = 32'h0;  // 32'h0742e5eb;
    ram_cell[      69] = 32'h0;  // 32'h0b333a65;
    ram_cell[      70] = 32'h0;  // 32'h8a747299;
    ram_cell[      71] = 32'h0;  // 32'h2dbe6c8d;
    ram_cell[      72] = 32'h0;  // 32'h54e5888a;
    ram_cell[      73] = 32'h0;  // 32'hbd611d4f;
    ram_cell[      74] = 32'h0;  // 32'hf66dbb80;
    ram_cell[      75] = 32'h0;  // 32'h9da0ffa4;
    ram_cell[      76] = 32'h0;  // 32'h2911fe60;
    ram_cell[      77] = 32'h0;  // 32'h8e79268a;
    ram_cell[      78] = 32'h0;  // 32'he9e07a73;
    ram_cell[      79] = 32'h0;  // 32'h64ac168d;
    ram_cell[      80] = 32'h0;  // 32'h188ce858;
    ram_cell[      81] = 32'h0;  // 32'ha089737f;
    ram_cell[      82] = 32'h0;  // 32'h8d5890e2;
    ram_cell[      83] = 32'h0;  // 32'h5b2bc019;
    ram_cell[      84] = 32'h0;  // 32'hd09de5d3;
    ram_cell[      85] = 32'h0;  // 32'h61150c97;
    ram_cell[      86] = 32'h0;  // 32'hbd24e997;
    ram_cell[      87] = 32'h0;  // 32'h0bb91b29;
    ram_cell[      88] = 32'h0;  // 32'h39e0c0d7;
    ram_cell[      89] = 32'h0;  // 32'h370775fb;
    ram_cell[      90] = 32'h0;  // 32'h23e567e0;
    ram_cell[      91] = 32'h0;  // 32'h636788b4;
    ram_cell[      92] = 32'h0;  // 32'h5bfb48bf;
    ram_cell[      93] = 32'h0;  // 32'hf746a6de;
    ram_cell[      94] = 32'h0;  // 32'hed4ad7f1;
    ram_cell[      95] = 32'h0;  // 32'h67f35fde;
    ram_cell[      96] = 32'h0;  // 32'h82001b56;
    ram_cell[      97] = 32'h0;  // 32'h58d3a032;
    ram_cell[      98] = 32'h0;  // 32'h75e9cf29;
    ram_cell[      99] = 32'h0;  // 32'h3644e671;
    ram_cell[     100] = 32'h0;  // 32'h078566c9;
    ram_cell[     101] = 32'h0;  // 32'hc4a22142;
    ram_cell[     102] = 32'h0;  // 32'h46ade047;
    ram_cell[     103] = 32'h0;  // 32'hf593c183;
    ram_cell[     104] = 32'h0;  // 32'h4a02c526;
    ram_cell[     105] = 32'h0;  // 32'h429e2c72;
    ram_cell[     106] = 32'h0;  // 32'h2103d070;
    ram_cell[     107] = 32'h0;  // 32'hc5cec9a0;
    ram_cell[     108] = 32'h0;  // 32'hfda80392;
    ram_cell[     109] = 32'h0;  // 32'he45eeed5;
    ram_cell[     110] = 32'h0;  // 32'hb19b564d;
    ram_cell[     111] = 32'h0;  // 32'hc2d24811;
    ram_cell[     112] = 32'h0;  // 32'h7dfa1f86;
    ram_cell[     113] = 32'h0;  // 32'h6c6113df;
    ram_cell[     114] = 32'h0;  // 32'h59f8fc1f;
    ram_cell[     115] = 32'h0;  // 32'h08f0dec8;
    ram_cell[     116] = 32'h0;  // 32'h30840770;
    ram_cell[     117] = 32'h0;  // 32'hd801cbf9;
    ram_cell[     118] = 32'h0;  // 32'hf980ca46;
    ram_cell[     119] = 32'h0;  // 32'h93cbfa10;
    ram_cell[     120] = 32'h0;  // 32'h148ad439;
    ram_cell[     121] = 32'h0;  // 32'hc2095e08;
    ram_cell[     122] = 32'h0;  // 32'hd6b2579a;
    ram_cell[     123] = 32'h0;  // 32'hc12e5360;
    ram_cell[     124] = 32'h0;  // 32'ha10d38ab;
    ram_cell[     125] = 32'h0;  // 32'h34ce0e89;
    ram_cell[     126] = 32'h0;  // 32'h38a75320;
    ram_cell[     127] = 32'h0;  // 32'h39c704ed;
    ram_cell[     128] = 32'h0;  // 32'h475b9efb;
    ram_cell[     129] = 32'h0;  // 32'h2a19f11f;
    ram_cell[     130] = 32'h0;  // 32'hdcb44729;
    ram_cell[     131] = 32'h0;  // 32'h39f25153;
    ram_cell[     132] = 32'h0;  // 32'hd4c9074b;
    ram_cell[     133] = 32'h0;  // 32'hbb28497b;
    ram_cell[     134] = 32'h0;  // 32'he6da0637;
    ram_cell[     135] = 32'h0;  // 32'h17fda05f;
    ram_cell[     136] = 32'h0;  // 32'h6c8e9136;
    ram_cell[     137] = 32'h0;  // 32'hf65fd9bc;
    ram_cell[     138] = 32'h0;  // 32'h820da878;
    ram_cell[     139] = 32'h0;  // 32'h337800c8;
    ram_cell[     140] = 32'h0;  // 32'h992a1f40;
    ram_cell[     141] = 32'h0;  // 32'h1d36bc3d;
    ram_cell[     142] = 32'h0;  // 32'h985b8d2a;
    ram_cell[     143] = 32'h0;  // 32'h852d5b07;
    ram_cell[     144] = 32'h0;  // 32'h8fc79336;
    ram_cell[     145] = 32'h0;  // 32'hd2cb795a;
    ram_cell[     146] = 32'h0;  // 32'h0033ddba;
    ram_cell[     147] = 32'h0;  // 32'h107b5e31;
    ram_cell[     148] = 32'h0;  // 32'h2141205e;
    ram_cell[     149] = 32'h0;  // 32'he49d06d6;
    ram_cell[     150] = 32'h0;  // 32'h23da9c63;
    ram_cell[     151] = 32'h0;  // 32'hc51fc5fb;
    ram_cell[     152] = 32'h0;  // 32'hc63c07ed;
    ram_cell[     153] = 32'h0;  // 32'h8faed34c;
    ram_cell[     154] = 32'h0;  // 32'h7fd65b51;
    ram_cell[     155] = 32'h0;  // 32'he8a73a27;
    ram_cell[     156] = 32'h0;  // 32'h82da2c7b;
    ram_cell[     157] = 32'h0;  // 32'h458ca77e;
    ram_cell[     158] = 32'h0;  // 32'h02116332;
    ram_cell[     159] = 32'h0;  // 32'h64896303;
    ram_cell[     160] = 32'h0;  // 32'h2a9e85b3;
    ram_cell[     161] = 32'h0;  // 32'h70e4c706;
    ram_cell[     162] = 32'h0;  // 32'hd49db4f4;
    ram_cell[     163] = 32'h0;  // 32'h26bb176a;
    ram_cell[     164] = 32'h0;  // 32'h0bd39a75;
    ram_cell[     165] = 32'h0;  // 32'h454f2607;
    ram_cell[     166] = 32'h0;  // 32'h2601bc6a;
    ram_cell[     167] = 32'h0;  // 32'h444cfb6c;
    ram_cell[     168] = 32'h0;  // 32'h3fed62f4;
    ram_cell[     169] = 32'h0;  // 32'ha74c732d;
    ram_cell[     170] = 32'h0;  // 32'h26bbcc1c;
    ram_cell[     171] = 32'h0;  // 32'hd3287f70;
    ram_cell[     172] = 32'h0;  // 32'h064d840e;
    ram_cell[     173] = 32'h0;  // 32'h03056864;
    ram_cell[     174] = 32'h0;  // 32'h0c5e12ed;
    ram_cell[     175] = 32'h0;  // 32'h1746cbb5;
    ram_cell[     176] = 32'h0;  // 32'h7f39e502;
    ram_cell[     177] = 32'h0;  // 32'hd82bcece;
    ram_cell[     178] = 32'h0;  // 32'h99243c74;
    ram_cell[     179] = 32'h0;  // 32'h83d01aa8;
    ram_cell[     180] = 32'h0;  // 32'h4f0a85dd;
    ram_cell[     181] = 32'h0;  // 32'h2c77d5ff;
    ram_cell[     182] = 32'h0;  // 32'h51fb889f;
    ram_cell[     183] = 32'h0;  // 32'hbcd5413a;
    ram_cell[     184] = 32'h0;  // 32'h64e27e1b;
    ram_cell[     185] = 32'h0;  // 32'h945beec8;
    ram_cell[     186] = 32'h0;  // 32'h63bf3c94;
    ram_cell[     187] = 32'h0;  // 32'hbc219170;
    ram_cell[     188] = 32'h0;  // 32'h6e4369a4;
    ram_cell[     189] = 32'h0;  // 32'h84cbcf0b;
    ram_cell[     190] = 32'h0;  // 32'h50d17614;
    ram_cell[     191] = 32'h0;  // 32'h833bc41e;
    ram_cell[     192] = 32'h0;  // 32'h78b4b928;
    ram_cell[     193] = 32'h0;  // 32'h4a70ab1b;
    ram_cell[     194] = 32'h0;  // 32'h9c874346;
    ram_cell[     195] = 32'h0;  // 32'h9cf8c326;
    ram_cell[     196] = 32'h0;  // 32'h4a4d24c5;
    ram_cell[     197] = 32'h0;  // 32'hcfce7050;
    ram_cell[     198] = 32'h0;  // 32'h17902d25;
    ram_cell[     199] = 32'h0;  // 32'h015b5ffa;
    ram_cell[     200] = 32'h0;  // 32'hc016f091;
    ram_cell[     201] = 32'h0;  // 32'h0aa89bb4;
    ram_cell[     202] = 32'h0;  // 32'h6726a04d;
    ram_cell[     203] = 32'h0;  // 32'h1c123f48;
    ram_cell[     204] = 32'h0;  // 32'h002a5742;
    ram_cell[     205] = 32'h0;  // 32'ha1003747;
    ram_cell[     206] = 32'h0;  // 32'hf31dc84d;
    ram_cell[     207] = 32'h0;  // 32'h1f6fdb93;
    ram_cell[     208] = 32'h0;  // 32'h61f14182;
    ram_cell[     209] = 32'h0;  // 32'h124f5150;
    ram_cell[     210] = 32'h0;  // 32'he8aac64b;
    ram_cell[     211] = 32'h0;  // 32'hb5ad6d83;
    ram_cell[     212] = 32'h0;  // 32'h13e7f80e;
    ram_cell[     213] = 32'h0;  // 32'hb4074451;
    ram_cell[     214] = 32'h0;  // 32'hb46a24b6;
    ram_cell[     215] = 32'h0;  // 32'h1ceb0a88;
    ram_cell[     216] = 32'h0;  // 32'h7c632fd6;
    ram_cell[     217] = 32'h0;  // 32'h556807ba;
    ram_cell[     218] = 32'h0;  // 32'h94f051e8;
    ram_cell[     219] = 32'h0;  // 32'h66819167;
    ram_cell[     220] = 32'h0;  // 32'h9fabbaee;
    ram_cell[     221] = 32'h0;  // 32'h09edd1dd;
    ram_cell[     222] = 32'h0;  // 32'he614dbe9;
    ram_cell[     223] = 32'h0;  // 32'hb7aa8163;
    ram_cell[     224] = 32'h0;  // 32'hc2b0d271;
    ram_cell[     225] = 32'h0;  // 32'hcb73c71a;
    ram_cell[     226] = 32'h0;  // 32'h9b500085;
    ram_cell[     227] = 32'h0;  // 32'hcbceda2b;
    ram_cell[     228] = 32'h0;  // 32'hc842d4bd;
    ram_cell[     229] = 32'h0;  // 32'h48860367;
    ram_cell[     230] = 32'h0;  // 32'hd0b7e0e1;
    ram_cell[     231] = 32'h0;  // 32'h0ce6c20a;
    ram_cell[     232] = 32'h0;  // 32'h37308527;
    ram_cell[     233] = 32'h0;  // 32'hd4818059;
    ram_cell[     234] = 32'h0;  // 32'hadbc1747;
    ram_cell[     235] = 32'h0;  // 32'h36625f0a;
    ram_cell[     236] = 32'h0;  // 32'h03af7b59;
    ram_cell[     237] = 32'h0;  // 32'hb3403a86;
    ram_cell[     238] = 32'h0;  // 32'h2311229d;
    ram_cell[     239] = 32'h0;  // 32'ha2598ffb;
    ram_cell[     240] = 32'h0;  // 32'h86eed1ba;
    ram_cell[     241] = 32'h0;  // 32'hf4f77ae9;
    ram_cell[     242] = 32'h0;  // 32'h796064e4;
    ram_cell[     243] = 32'h0;  // 32'h60fb3a31;
    ram_cell[     244] = 32'h0;  // 32'hbccc87b3;
    ram_cell[     245] = 32'h0;  // 32'h3e0558c6;
    ram_cell[     246] = 32'h0;  // 32'he583e84b;
    ram_cell[     247] = 32'h0;  // 32'h7e68e7c8;
    ram_cell[     248] = 32'h0;  // 32'h28529915;
    ram_cell[     249] = 32'h0;  // 32'h662b08a9;
    ram_cell[     250] = 32'h0;  // 32'hcff18716;
    ram_cell[     251] = 32'h0;  // 32'h57835f50;
    ram_cell[     252] = 32'h0;  // 32'h3611820d;
    ram_cell[     253] = 32'h0;  // 32'hccaf02a4;
    ram_cell[     254] = 32'h0;  // 32'h7bda3293;
    ram_cell[     255] = 32'h0;  // 32'h710a9013;
    // src matrix A
    ram_cell[     256] = 32'h040324f7;
    ram_cell[     257] = 32'h95ba51b9;
    ram_cell[     258] = 32'h95e2eb8b;
    ram_cell[     259] = 32'h5e53247b;
    ram_cell[     260] = 32'h3e3b092f;
    ram_cell[     261] = 32'h061b4711;
    ram_cell[     262] = 32'h941a155e;
    ram_cell[     263] = 32'hac791354;
    ram_cell[     264] = 32'ha4ee8ca4;
    ram_cell[     265] = 32'h82c28517;
    ram_cell[     266] = 32'hc49d5659;
    ram_cell[     267] = 32'h30aad2ba;
    ram_cell[     268] = 32'h8ed66066;
    ram_cell[     269] = 32'h51e5affc;
    ram_cell[     270] = 32'h5e3c78cd;
    ram_cell[     271] = 32'hcd35fc79;
    ram_cell[     272] = 32'h43291236;
    ram_cell[     273] = 32'hbd6244ea;
    ram_cell[     274] = 32'hb486f3ea;
    ram_cell[     275] = 32'h447473eb;
    ram_cell[     276] = 32'h45890fce;
    ram_cell[     277] = 32'h8a8c589c;
    ram_cell[     278] = 32'h14eaabee;
    ram_cell[     279] = 32'h4e7e9edb;
    ram_cell[     280] = 32'h32e102c4;
    ram_cell[     281] = 32'h08cda4bb;
    ram_cell[     282] = 32'h486deea4;
    ram_cell[     283] = 32'h67991139;
    ram_cell[     284] = 32'hca57f793;
    ram_cell[     285] = 32'h4e81edc6;
    ram_cell[     286] = 32'hd821c107;
    ram_cell[     287] = 32'h3c715fd8;
    ram_cell[     288] = 32'hdec840fd;
    ram_cell[     289] = 32'h73e80242;
    ram_cell[     290] = 32'ha0f11455;
    ram_cell[     291] = 32'h975147bb;
    ram_cell[     292] = 32'h5573db67;
    ram_cell[     293] = 32'h2f04b2dc;
    ram_cell[     294] = 32'h635b926c;
    ram_cell[     295] = 32'hd58d6dc5;
    ram_cell[     296] = 32'ha8623473;
    ram_cell[     297] = 32'h847e30e7;
    ram_cell[     298] = 32'hf79ed5c9;
    ram_cell[     299] = 32'h264f60b4;
    ram_cell[     300] = 32'h232ec952;
    ram_cell[     301] = 32'had85543a;
    ram_cell[     302] = 32'h297f6f9d;
    ram_cell[     303] = 32'hda825908;
    ram_cell[     304] = 32'hc9f2cd83;
    ram_cell[     305] = 32'h9fdd7fd1;
    ram_cell[     306] = 32'hb860a37a;
    ram_cell[     307] = 32'h5ff92faa;
    ram_cell[     308] = 32'hd78ecb91;
    ram_cell[     309] = 32'h07c4e7b2;
    ram_cell[     310] = 32'h2ca9abb0;
    ram_cell[     311] = 32'h49d41abb;
    ram_cell[     312] = 32'h2e15b048;
    ram_cell[     313] = 32'h37fa8cea;
    ram_cell[     314] = 32'hb17493c2;
    ram_cell[     315] = 32'hbb59260d;
    ram_cell[     316] = 32'h3721cf6d;
    ram_cell[     317] = 32'h0ebfbc6e;
    ram_cell[     318] = 32'h0b23ecaf;
    ram_cell[     319] = 32'h4aec9398;
    ram_cell[     320] = 32'h5b080103;
    ram_cell[     321] = 32'h7134489f;
    ram_cell[     322] = 32'h3eb69712;
    ram_cell[     323] = 32'h1a7cd4d3;
    ram_cell[     324] = 32'h1ad59280;
    ram_cell[     325] = 32'hb9e33e81;
    ram_cell[     326] = 32'h04d8635e;
    ram_cell[     327] = 32'h743d55c9;
    ram_cell[     328] = 32'h9b1a8daa;
    ram_cell[     329] = 32'hbef51b46;
    ram_cell[     330] = 32'h5177dd87;
    ram_cell[     331] = 32'h5285e853;
    ram_cell[     332] = 32'h8ef96f1c;
    ram_cell[     333] = 32'h639e10ac;
    ram_cell[     334] = 32'h0ba4c748;
    ram_cell[     335] = 32'h688f7434;
    ram_cell[     336] = 32'h7412991b;
    ram_cell[     337] = 32'h4f818e7f;
    ram_cell[     338] = 32'he90961d1;
    ram_cell[     339] = 32'hf9adc517;
    ram_cell[     340] = 32'h1744c6f3;
    ram_cell[     341] = 32'h5a025f5f;
    ram_cell[     342] = 32'h9d8b6558;
    ram_cell[     343] = 32'hb24856c0;
    ram_cell[     344] = 32'h0d52e4e4;
    ram_cell[     345] = 32'hb10f0438;
    ram_cell[     346] = 32'hd9d9858b;
    ram_cell[     347] = 32'ha4a7939a;
    ram_cell[     348] = 32'hf2810850;
    ram_cell[     349] = 32'h5f86c4ff;
    ram_cell[     350] = 32'hd1852e38;
    ram_cell[     351] = 32'hacd8f2e9;
    ram_cell[     352] = 32'h240bcd5e;
    ram_cell[     353] = 32'he7e8574a;
    ram_cell[     354] = 32'hc60adf2a;
    ram_cell[     355] = 32'hca678dd1;
    ram_cell[     356] = 32'h7cdecd7b;
    ram_cell[     357] = 32'hbc6f0dd7;
    ram_cell[     358] = 32'hd2e73bb3;
    ram_cell[     359] = 32'he8a3f6a6;
    ram_cell[     360] = 32'hc8487854;
    ram_cell[     361] = 32'hecd9cd45;
    ram_cell[     362] = 32'he6fbd002;
    ram_cell[     363] = 32'h08121236;
    ram_cell[     364] = 32'h71885294;
    ram_cell[     365] = 32'hf419b52f;
    ram_cell[     366] = 32'h04630d50;
    ram_cell[     367] = 32'hb4627045;
    ram_cell[     368] = 32'hb5fa96f9;
    ram_cell[     369] = 32'he2e4e4aa;
    ram_cell[     370] = 32'hf377e909;
    ram_cell[     371] = 32'h8b7ef235;
    ram_cell[     372] = 32'h79f89a25;
    ram_cell[     373] = 32'h8c836b1d;
    ram_cell[     374] = 32'h468ce94a;
    ram_cell[     375] = 32'h1a979733;
    ram_cell[     376] = 32'hbae6f0ec;
    ram_cell[     377] = 32'ha0508cc9;
    ram_cell[     378] = 32'h55ea2cbe;
    ram_cell[     379] = 32'hb4ac8d4c;
    ram_cell[     380] = 32'h5a1d25a2;
    ram_cell[     381] = 32'h97893a0e;
    ram_cell[     382] = 32'ha8f1cf38;
    ram_cell[     383] = 32'hd098c959;
    ram_cell[     384] = 32'hd45df87d;
    ram_cell[     385] = 32'h21cb9a32;
    ram_cell[     386] = 32'h462f6526;
    ram_cell[     387] = 32'h1fe3d3ba;
    ram_cell[     388] = 32'h8fab24f4;
    ram_cell[     389] = 32'hfa07ae9d;
    ram_cell[     390] = 32'ha1d2baf9;
    ram_cell[     391] = 32'h53c0a40a;
    ram_cell[     392] = 32'h21837d92;
    ram_cell[     393] = 32'hde1dc35a;
    ram_cell[     394] = 32'hcec85dfb;
    ram_cell[     395] = 32'hfda54081;
    ram_cell[     396] = 32'h5e9ebaa2;
    ram_cell[     397] = 32'h76007ac0;
    ram_cell[     398] = 32'h2317d0db;
    ram_cell[     399] = 32'hd734db3e;
    ram_cell[     400] = 32'hd8d9c0e0;
    ram_cell[     401] = 32'hb1bd74bf;
    ram_cell[     402] = 32'h6c5524aa;
    ram_cell[     403] = 32'h4ac19a1e;
    ram_cell[     404] = 32'h0ce92679;
    ram_cell[     405] = 32'hf57eb997;
    ram_cell[     406] = 32'haa59c8e0;
    ram_cell[     407] = 32'h281816f5;
    ram_cell[     408] = 32'ha326358d;
    ram_cell[     409] = 32'h0048543d;
    ram_cell[     410] = 32'h7fdd4e5c;
    ram_cell[     411] = 32'he7d16969;
    ram_cell[     412] = 32'h761ffb81;
    ram_cell[     413] = 32'h3ae0f260;
    ram_cell[     414] = 32'haa6ebc4c;
    ram_cell[     415] = 32'h52c57bf4;
    ram_cell[     416] = 32'h1b289d85;
    ram_cell[     417] = 32'h7d03c131;
    ram_cell[     418] = 32'h3651ca83;
    ram_cell[     419] = 32'ha87587a1;
    ram_cell[     420] = 32'h5ef7490e;
    ram_cell[     421] = 32'h9dcd91d6;
    ram_cell[     422] = 32'h7bf79ba6;
    ram_cell[     423] = 32'h01f3695d;
    ram_cell[     424] = 32'h18f5603d;
    ram_cell[     425] = 32'h761db965;
    ram_cell[     426] = 32'hcedaff7f;
    ram_cell[     427] = 32'h233ea125;
    ram_cell[     428] = 32'he53f8fa5;
    ram_cell[     429] = 32'h7cf84a65;
    ram_cell[     430] = 32'h8e964a2a;
    ram_cell[     431] = 32'h9347ad9e;
    ram_cell[     432] = 32'he588dc84;
    ram_cell[     433] = 32'h610d9138;
    ram_cell[     434] = 32'h82cb1071;
    ram_cell[     435] = 32'he21d15c9;
    ram_cell[     436] = 32'hc82a9971;
    ram_cell[     437] = 32'h96cfbcba;
    ram_cell[     438] = 32'hfcc590a4;
    ram_cell[     439] = 32'h38cdf6ee;
    ram_cell[     440] = 32'hd0e02cd7;
    ram_cell[     441] = 32'h0df830bb;
    ram_cell[     442] = 32'h95a8013d;
    ram_cell[     443] = 32'hd2b62c58;
    ram_cell[     444] = 32'hf4a25fb0;
    ram_cell[     445] = 32'h83eafa5a;
    ram_cell[     446] = 32'h4320c99c;
    ram_cell[     447] = 32'hda190df4;
    ram_cell[     448] = 32'h6a469c8c;
    ram_cell[     449] = 32'h082749ed;
    ram_cell[     450] = 32'h43e1ea8d;
    ram_cell[     451] = 32'had42ae80;
    ram_cell[     452] = 32'h5a1ff934;
    ram_cell[     453] = 32'h30d26038;
    ram_cell[     454] = 32'ha688d3b5;
    ram_cell[     455] = 32'h53a25522;
    ram_cell[     456] = 32'hc5d86a56;
    ram_cell[     457] = 32'h26082314;
    ram_cell[     458] = 32'h78e242ec;
    ram_cell[     459] = 32'h032046f6;
    ram_cell[     460] = 32'h2b284752;
    ram_cell[     461] = 32'h0b76f812;
    ram_cell[     462] = 32'h13c7708e;
    ram_cell[     463] = 32'hf5f068a0;
    ram_cell[     464] = 32'h8b1c548b;
    ram_cell[     465] = 32'h5df33e74;
    ram_cell[     466] = 32'h52424c05;
    ram_cell[     467] = 32'hc64de97b;
    ram_cell[     468] = 32'h92fef875;
    ram_cell[     469] = 32'hdb397d1f;
    ram_cell[     470] = 32'h67b85127;
    ram_cell[     471] = 32'h7184f26a;
    ram_cell[     472] = 32'h07e1f6f4;
    ram_cell[     473] = 32'h3755e752;
    ram_cell[     474] = 32'h467f18d5;
    ram_cell[     475] = 32'hbb681ea7;
    ram_cell[     476] = 32'h4af8cca3;
    ram_cell[     477] = 32'h68418a35;
    ram_cell[     478] = 32'h77691c71;
    ram_cell[     479] = 32'h6a310833;
    ram_cell[     480] = 32'h8fc3db53;
    ram_cell[     481] = 32'h362707aa;
    ram_cell[     482] = 32'h311c2d3f;
    ram_cell[     483] = 32'h96e0c8ac;
    ram_cell[     484] = 32'h8e5e728e;
    ram_cell[     485] = 32'h59fabc2b;
    ram_cell[     486] = 32'h2fc91cc3;
    ram_cell[     487] = 32'hc6eac24d;
    ram_cell[     488] = 32'h4749f07a;
    ram_cell[     489] = 32'hfc6a19e4;
    ram_cell[     490] = 32'h4f06c1b4;
    ram_cell[     491] = 32'h5f7cd7b3;
    ram_cell[     492] = 32'h75459c9f;
    ram_cell[     493] = 32'h24f20d44;
    ram_cell[     494] = 32'h6aedb9f4;
    ram_cell[     495] = 32'h5f322fa0;
    ram_cell[     496] = 32'h3dcc9b9f;
    ram_cell[     497] = 32'h64595772;
    ram_cell[     498] = 32'hddab5b69;
    ram_cell[     499] = 32'he86b2818;
    ram_cell[     500] = 32'hf70014ed;
    ram_cell[     501] = 32'h030e11ab;
    ram_cell[     502] = 32'h55ff4354;
    ram_cell[     503] = 32'h2a13beea;
    ram_cell[     504] = 32'h03817e00;
    ram_cell[     505] = 32'h131e858b;
    ram_cell[     506] = 32'hacb73b5a;
    ram_cell[     507] = 32'hccfb8dd3;
    ram_cell[     508] = 32'he36a92f0;
    ram_cell[     509] = 32'hde08d9f0;
    ram_cell[     510] = 32'h2e8b13ab;
    ram_cell[     511] = 32'h24068649;
    // src matrix B
    ram_cell[     512] = 32'h2213b392;
    ram_cell[     513] = 32'hc7deca0c;
    ram_cell[     514] = 32'h0eb6b9f2;
    ram_cell[     515] = 32'h06699750;
    ram_cell[     516] = 32'hd4e2644f;
    ram_cell[     517] = 32'hb15562e0;
    ram_cell[     518] = 32'h42943992;
    ram_cell[     519] = 32'h5b6dc9e7;
    ram_cell[     520] = 32'hc7b7d5ea;
    ram_cell[     521] = 32'h2181df84;
    ram_cell[     522] = 32'h9b9ec9fb;
    ram_cell[     523] = 32'hb0ed9225;
    ram_cell[     524] = 32'h7ee49910;
    ram_cell[     525] = 32'haba6937b;
    ram_cell[     526] = 32'hcaa65d0d;
    ram_cell[     527] = 32'h948839aa;
    ram_cell[     528] = 32'hdaab165a;
    ram_cell[     529] = 32'h62e2ce25;
    ram_cell[     530] = 32'hb1935b42;
    ram_cell[     531] = 32'hb9fa04d3;
    ram_cell[     532] = 32'h3ebb7d70;
    ram_cell[     533] = 32'h3b4f8a1f;
    ram_cell[     534] = 32'h50848a52;
    ram_cell[     535] = 32'hc4e2a2d1;
    ram_cell[     536] = 32'h7c6d0a8c;
    ram_cell[     537] = 32'h4b0d6c5f;
    ram_cell[     538] = 32'haf754ba5;
    ram_cell[     539] = 32'h18cb65f3;
    ram_cell[     540] = 32'h50732ede;
    ram_cell[     541] = 32'h966a69f9;
    ram_cell[     542] = 32'h6b44e381;
    ram_cell[     543] = 32'hbcc093c8;
    ram_cell[     544] = 32'hff9dc5de;
    ram_cell[     545] = 32'hcd386e1f;
    ram_cell[     546] = 32'h58543f28;
    ram_cell[     547] = 32'h5c3b7b94;
    ram_cell[     548] = 32'hcdc23516;
    ram_cell[     549] = 32'hdba726f7;
    ram_cell[     550] = 32'h33c31466;
    ram_cell[     551] = 32'h7b33f821;
    ram_cell[     552] = 32'h08534ab9;
    ram_cell[     553] = 32'h454011c7;
    ram_cell[     554] = 32'hb853224d;
    ram_cell[     555] = 32'h62403584;
    ram_cell[     556] = 32'h0a8417b4;
    ram_cell[     557] = 32'h5d03df4e;
    ram_cell[     558] = 32'h317032e3;
    ram_cell[     559] = 32'h1eb3f356;
    ram_cell[     560] = 32'hbd968866;
    ram_cell[     561] = 32'hefe9c6fa;
    ram_cell[     562] = 32'h7fed0bba;
    ram_cell[     563] = 32'h5240159c;
    ram_cell[     564] = 32'h89ba5f3d;
    ram_cell[     565] = 32'h35d8c6c1;
    ram_cell[     566] = 32'h965478cd;
    ram_cell[     567] = 32'haf9da6a8;
    ram_cell[     568] = 32'hd8d1a138;
    ram_cell[     569] = 32'h003ba907;
    ram_cell[     570] = 32'h999ef979;
    ram_cell[     571] = 32'h7f47e1a3;
    ram_cell[     572] = 32'h33ff6865;
    ram_cell[     573] = 32'hd6fbb0a2;
    ram_cell[     574] = 32'hc202306c;
    ram_cell[     575] = 32'h6cf70cae;
    ram_cell[     576] = 32'h5e88e052;
    ram_cell[     577] = 32'h08cf2dce;
    ram_cell[     578] = 32'h1d525cf4;
    ram_cell[     579] = 32'hd5c583a8;
    ram_cell[     580] = 32'h3303709f;
    ram_cell[     581] = 32'hef46d0c8;
    ram_cell[     582] = 32'hd443a2fe;
    ram_cell[     583] = 32'h1e1935d8;
    ram_cell[     584] = 32'h5bb0d854;
    ram_cell[     585] = 32'h734a2042;
    ram_cell[     586] = 32'h24ea0a52;
    ram_cell[     587] = 32'h1fe6819a;
    ram_cell[     588] = 32'h9c099baa;
    ram_cell[     589] = 32'ha3a225a1;
    ram_cell[     590] = 32'h2d1c2b44;
    ram_cell[     591] = 32'ha2800ff3;
    ram_cell[     592] = 32'hf089115e;
    ram_cell[     593] = 32'h9a02254b;
    ram_cell[     594] = 32'h0e5cc816;
    ram_cell[     595] = 32'h155c965d;
    ram_cell[     596] = 32'hf576c34b;
    ram_cell[     597] = 32'heb3782ef;
    ram_cell[     598] = 32'h78ecb3dc;
    ram_cell[     599] = 32'h69141b79;
    ram_cell[     600] = 32'h931db207;
    ram_cell[     601] = 32'h63dd0037;
    ram_cell[     602] = 32'ha4fd7c0b;
    ram_cell[     603] = 32'h18d13146;
    ram_cell[     604] = 32'h8e4793eb;
    ram_cell[     605] = 32'h17d61675;
    ram_cell[     606] = 32'hb91d4559;
    ram_cell[     607] = 32'h6aa6d49f;
    ram_cell[     608] = 32'h96690b76;
    ram_cell[     609] = 32'he7bec153;
    ram_cell[     610] = 32'hc5ba09f6;
    ram_cell[     611] = 32'h717afd83;
    ram_cell[     612] = 32'h756d06a5;
    ram_cell[     613] = 32'hfa31e280;
    ram_cell[     614] = 32'h83de9e4f;
    ram_cell[     615] = 32'h71947f62;
    ram_cell[     616] = 32'h2a05b57c;
    ram_cell[     617] = 32'he5f66e98;
    ram_cell[     618] = 32'hc9c5d0df;
    ram_cell[     619] = 32'h24ae4f2d;
    ram_cell[     620] = 32'ha07273dc;
    ram_cell[     621] = 32'h34b73222;
    ram_cell[     622] = 32'hc92a6223;
    ram_cell[     623] = 32'h18ab4f0d;
    ram_cell[     624] = 32'h16d8f280;
    ram_cell[     625] = 32'h1b4e933f;
    ram_cell[     626] = 32'h5dbc34cd;
    ram_cell[     627] = 32'h13f30f92;
    ram_cell[     628] = 32'h05405229;
    ram_cell[     629] = 32'h148070ca;
    ram_cell[     630] = 32'h56805eb5;
    ram_cell[     631] = 32'h2c81fdb4;
    ram_cell[     632] = 32'h05ff38e4;
    ram_cell[     633] = 32'h4a0b530a;
    ram_cell[     634] = 32'h3b0ef864;
    ram_cell[     635] = 32'ha2782d7c;
    ram_cell[     636] = 32'h6ea1c17d;
    ram_cell[     637] = 32'h8b571d41;
    ram_cell[     638] = 32'h18546df6;
    ram_cell[     639] = 32'h0cf8ee9e;
    ram_cell[     640] = 32'hc0e7226c;
    ram_cell[     641] = 32'h9febdcf9;
    ram_cell[     642] = 32'h7ee9dfb5;
    ram_cell[     643] = 32'hf8bf787c;
    ram_cell[     644] = 32'h05d86d3f;
    ram_cell[     645] = 32'h8a2c4eb4;
    ram_cell[     646] = 32'hc310a29b;
    ram_cell[     647] = 32'h3d14e82c;
    ram_cell[     648] = 32'hb664c58a;
    ram_cell[     649] = 32'hcd74b56f;
    ram_cell[     650] = 32'hfff128aa;
    ram_cell[     651] = 32'he1bf9e26;
    ram_cell[     652] = 32'hb5a8bce0;
    ram_cell[     653] = 32'h4fd537c7;
    ram_cell[     654] = 32'hb3b36411;
    ram_cell[     655] = 32'h06abd2e3;
    ram_cell[     656] = 32'h2b51c54d;
    ram_cell[     657] = 32'h8a1ed298;
    ram_cell[     658] = 32'h901d36a8;
    ram_cell[     659] = 32'h70375470;
    ram_cell[     660] = 32'h702b0f53;
    ram_cell[     661] = 32'h00e5ea25;
    ram_cell[     662] = 32'hf83bfd88;
    ram_cell[     663] = 32'hab6b8582;
    ram_cell[     664] = 32'h2226ad1f;
    ram_cell[     665] = 32'ha436f2e4;
    ram_cell[     666] = 32'h8a9f0d92;
    ram_cell[     667] = 32'h638e7dbe;
    ram_cell[     668] = 32'h337b2758;
    ram_cell[     669] = 32'h88fbe41e;
    ram_cell[     670] = 32'h54c87cbc;
    ram_cell[     671] = 32'h2b7540ff;
    ram_cell[     672] = 32'h5871d6ad;
    ram_cell[     673] = 32'h86cbb740;
    ram_cell[     674] = 32'h23d6b45f;
    ram_cell[     675] = 32'h6a330da8;
    ram_cell[     676] = 32'h2f9c663d;
    ram_cell[     677] = 32'hc1de78a6;
    ram_cell[     678] = 32'h69fe47ef;
    ram_cell[     679] = 32'ha285285d;
    ram_cell[     680] = 32'h29f4831f;
    ram_cell[     681] = 32'hcc0ad049;
    ram_cell[     682] = 32'h61f251a0;
    ram_cell[     683] = 32'hf89a07b5;
    ram_cell[     684] = 32'hf2880699;
    ram_cell[     685] = 32'h7cdee3a5;
    ram_cell[     686] = 32'hdec233b6;
    ram_cell[     687] = 32'h4d7a48a5;
    ram_cell[     688] = 32'hb56d43f3;
    ram_cell[     689] = 32'hc0c13fee;
    ram_cell[     690] = 32'ha107ead7;
    ram_cell[     691] = 32'h84386de6;
    ram_cell[     692] = 32'h897ed7f6;
    ram_cell[     693] = 32'hfd90ef80;
    ram_cell[     694] = 32'h8ccf889e;
    ram_cell[     695] = 32'h5f0c58c3;
    ram_cell[     696] = 32'h99f44470;
    ram_cell[     697] = 32'hc9e32033;
    ram_cell[     698] = 32'h5d05f37c;
    ram_cell[     699] = 32'ha91cab30;
    ram_cell[     700] = 32'h796e9b76;
    ram_cell[     701] = 32'h735fb7a1;
    ram_cell[     702] = 32'h5156a2de;
    ram_cell[     703] = 32'h3f08bc39;
    ram_cell[     704] = 32'h92a562fa;
    ram_cell[     705] = 32'h92b21300;
    ram_cell[     706] = 32'h7ec887f1;
    ram_cell[     707] = 32'h2b474997;
    ram_cell[     708] = 32'h1aa28921;
    ram_cell[     709] = 32'h15b150cf;
    ram_cell[     710] = 32'h1c2fd6ed;
    ram_cell[     711] = 32'h34faa4a8;
    ram_cell[     712] = 32'h56e29f57;
    ram_cell[     713] = 32'hb7eba752;
    ram_cell[     714] = 32'h0f5e8631;
    ram_cell[     715] = 32'hb9a2f2ac;
    ram_cell[     716] = 32'hcc8d552b;
    ram_cell[     717] = 32'hdc0bae1a;
    ram_cell[     718] = 32'hee5f416b;
    ram_cell[     719] = 32'h30a443ba;
    ram_cell[     720] = 32'hdccb4a16;
    ram_cell[     721] = 32'hba1d5510;
    ram_cell[     722] = 32'h27e67565;
    ram_cell[     723] = 32'h715372ee;
    ram_cell[     724] = 32'h946d616e;
    ram_cell[     725] = 32'h7b761130;
    ram_cell[     726] = 32'h73f700fb;
    ram_cell[     727] = 32'h6cef2ef3;
    ram_cell[     728] = 32'h9a89cce6;
    ram_cell[     729] = 32'hf5ea706b;
    ram_cell[     730] = 32'h65f9c579;
    ram_cell[     731] = 32'h7f0b8ff8;
    ram_cell[     732] = 32'h25de57ec;
    ram_cell[     733] = 32'h480fae44;
    ram_cell[     734] = 32'hcea30444;
    ram_cell[     735] = 32'haa660373;
    ram_cell[     736] = 32'h77961d8f;
    ram_cell[     737] = 32'hd1dc8ab9;
    ram_cell[     738] = 32'hdd49d381;
    ram_cell[     739] = 32'hf35f8b11;
    ram_cell[     740] = 32'hb57abebb;
    ram_cell[     741] = 32'h5e6e7e66;
    ram_cell[     742] = 32'h00f9372b;
    ram_cell[     743] = 32'h8f297989;
    ram_cell[     744] = 32'h0614b526;
    ram_cell[     745] = 32'h1c06e1c5;
    ram_cell[     746] = 32'h48de87c1;
    ram_cell[     747] = 32'h5d33effd;
    ram_cell[     748] = 32'hcf05d156;
    ram_cell[     749] = 32'h6103f2fb;
    ram_cell[     750] = 32'hb2477eb1;
    ram_cell[     751] = 32'h8ac81603;
    ram_cell[     752] = 32'he0db79b7;
    ram_cell[     753] = 32'ha9893c0a;
    ram_cell[     754] = 32'h9b3b1e48;
    ram_cell[     755] = 32'h37c609fb;
    ram_cell[     756] = 32'h6c8e27f2;
    ram_cell[     757] = 32'h49683e97;
    ram_cell[     758] = 32'ha963c6de;
    ram_cell[     759] = 32'hf7833c55;
    ram_cell[     760] = 32'h81462caa;
    ram_cell[     761] = 32'he3091219;
    ram_cell[     762] = 32'hea63899c;
    ram_cell[     763] = 32'h928d7e80;
    ram_cell[     764] = 32'h5381aaac;
    ram_cell[     765] = 32'hac91107d;
    ram_cell[     766] = 32'h33b215c7;
    ram_cell[     767] = 32'h27b22d6c;
end

endmodule

